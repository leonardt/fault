module myinv(
    input in_,
    output out
);

    assign out = ~in_;

endmodule
