module fatal_task;
    initial begin
        $fatal;
    end
endmodule
