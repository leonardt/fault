`timescale 1ns/1ns
module test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk_tb;

    reg [5:0] I [4:0][11:0][2:0];
    wire [5:0] O [4:0][11:0][2:0];

    

    test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk #(
        
    ) dut (
        .I(I),
        .O(O)
    );

    initial begin
        I[3][6][0] <= 6'd5;
        I[3][6][1] <= 6'd33;
        I[3][6][2] <= 6'd62;
        #1;
        if (!(O[3][6][0] === 6'd5)) begin
            $error("Failed on action=4 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][0].  Expected %x, got %x.", 6'd5, O[3][6][0]);
        end
        if (!(O[3][6][1] === 6'd33)) begin
            $error("Failed on action=5 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][1].  Expected %x, got %x.", 6'd33, O[3][6][1]);
        end
        if (!(O[3][6][2] === 6'd62)) begin
            $error("Failed on action=6 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][2].  Expected %x, got %x.", 6'd62, O[3][6][2]);
        end
        I[3][4][0] <= 6'd61;
        I[3][4][1] <= 6'd45;
        I[3][4][2] <= 6'd27;
        #1;
        if (!(O[3][4][0] === 6'd61)) begin
            $error("Failed on action=11 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][0].  Expected %x, got %x.", 6'd61, O[3][4][0]);
        end
        if (!(O[3][4][1] === 6'd45)) begin
            $error("Failed on action=12 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][1].  Expected %x, got %x.", 6'd45, O[3][4][1]);
        end
        if (!(O[3][4][2] === 6'd27)) begin
            $error("Failed on action=13 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][2].  Expected %x, got %x.", 6'd27, O[3][4][2]);
        end
        I[4][2][0] <= 6'd36;
        I[4][2][1] <= 6'd17;
        I[4][2][2] <= 6'd12;
        #1;
        if (!(O[4][2][0] === 6'd36)) begin
            $error("Failed on action=18 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][0].  Expected %x, got %x.", 6'd36, O[4][2][0]);
        end
        if (!(O[4][2][1] === 6'd17)) begin
            $error("Failed on action=19 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][1].  Expected %x, got %x.", 6'd17, O[4][2][1]);
        end
        if (!(O[4][2][2] === 6'd12)) begin
            $error("Failed on action=20 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][2].  Expected %x, got %x.", 6'd12, O[4][2][2]);
        end
        I[4][4][0] <= 6'd18;
        I[4][4][1] <= 6'd39;
        I[4][4][2] <= 6'd12;
        #1;
        if (!(O[4][4][0] === 6'd18)) begin
            $error("Failed on action=25 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][0].  Expected %x, got %x.", 6'd18, O[4][4][0]);
        end
        if (!(O[4][4][1] === 6'd39)) begin
            $error("Failed on action=26 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][1].  Expected %x, got %x.", 6'd39, O[4][4][1]);
        end
        if (!(O[4][4][2] === 6'd12)) begin
            $error("Failed on action=27 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][2].  Expected %x, got %x.", 6'd12, O[4][4][2]);
        end
        I[0][10][0] <= 6'd42;
        I[0][10][1] <= 6'd60;
        I[0][10][2] <= 6'd12;
        #1;
        if (!(O[0][10][0] === 6'd42)) begin
            $error("Failed on action=32 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][0].  Expected %x, got %x.", 6'd42, O[0][10][0]);
        end
        if (!(O[0][10][1] === 6'd60)) begin
            $error("Failed on action=33 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][1].  Expected %x, got %x.", 6'd60, O[0][10][1]);
        end
        if (!(O[0][10][2] === 6'd12)) begin
            $error("Failed on action=34 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][2].  Expected %x, got %x.", 6'd12, O[0][10][2]);
        end
        I[2][6][0] <= 6'd40;
        I[2][6][1] <= 6'd26;
        I[2][6][2] <= 6'd61;
        #1;
        if (!(O[2][6][0] === 6'd40)) begin
            $error("Failed on action=39 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][0].  Expected %x, got %x.", 6'd40, O[2][6][0]);
        end
        if (!(O[2][6][1] === 6'd26)) begin
            $error("Failed on action=40 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][1].  Expected %x, got %x.", 6'd26, O[2][6][1]);
        end
        if (!(O[2][6][2] === 6'd61)) begin
            $error("Failed on action=41 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][2].  Expected %x, got %x.", 6'd61, O[2][6][2]);
        end
        I[3][8][0] <= 6'd33;
        I[3][8][1] <= 6'd7;
        I[3][8][2] <= 6'd1;
        #1;
        if (!(O[3][8][0] === 6'd33)) begin
            $error("Failed on action=46 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][8][0].  Expected %x, got %x.", 6'd33, O[3][8][0]);
        end
        if (!(O[3][8][1] === 6'd7)) begin
            $error("Failed on action=47 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][8][1].  Expected %x, got %x.", 6'd7, O[3][8][1]);
        end
        if (!(O[3][8][2] === 6'd1)) begin
            $error("Failed on action=48 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][8][2].  Expected %x, got %x.", 6'd1, O[3][8][2]);
        end
        I[0][11][0] <= 6'd51;
        I[0][11][1] <= 6'd0;
        I[0][11][2] <= 6'd63;
        #1;
        if (!(O[0][11][0] === 6'd51)) begin
            $error("Failed on action=53 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][0].  Expected %x, got %x.", 6'd51, O[0][11][0]);
        end
        if (!(O[0][11][1] === 6'd0)) begin
            $error("Failed on action=54 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][1].  Expected %x, got %x.", 6'd0, O[0][11][1]);
        end
        if (!(O[0][11][2] === 6'd63)) begin
            $error("Failed on action=55 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][2].  Expected %x, got %x.", 6'd63, O[0][11][2]);
        end
        I[2][3][0] <= 6'd41;
        I[2][3][1] <= 6'd8;
        I[2][3][2] <= 6'd24;
        #1;
        if (!(O[2][3][0] === 6'd41)) begin
            $error("Failed on action=60 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][0].  Expected %x, got %x.", 6'd41, O[2][3][0]);
        end
        if (!(O[2][3][1] === 6'd8)) begin
            $error("Failed on action=61 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][1].  Expected %x, got %x.", 6'd8, O[2][3][1]);
        end
        if (!(O[2][3][2] === 6'd24)) begin
            $error("Failed on action=62 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][2].  Expected %x, got %x.", 6'd24, O[2][3][2]);
        end
        I[4][3][0] <= 6'd30;
        I[4][3][1] <= 6'd18;
        I[4][3][2] <= 6'd57;
        #1;
        if (!(O[4][3][0] === 6'd30)) begin
            $error("Failed on action=67 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][0].  Expected %x, got %x.", 6'd30, O[4][3][0]);
        end
        if (!(O[4][3][1] === 6'd18)) begin
            $error("Failed on action=68 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][1].  Expected %x, got %x.", 6'd18, O[4][3][1]);
        end
        if (!(O[4][3][2] === 6'd57)) begin
            $error("Failed on action=69 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][2].  Expected %x, got %x.", 6'd57, O[4][3][2]);
        end
        I[0][1][0] <= 6'd40;
        I[0][1][1] <= 6'd62;
        I[0][1][2] <= 6'd13;
        #1;
        if (!(O[0][1][0] === 6'd40)) begin
            $error("Failed on action=74 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][0].  Expected %x, got %x.", 6'd40, O[0][1][0]);
        end
        if (!(O[0][1][1] === 6'd62)) begin
            $error("Failed on action=75 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][1].  Expected %x, got %x.", 6'd62, O[0][1][1]);
        end
        if (!(O[0][1][2] === 6'd13)) begin
            $error("Failed on action=76 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][2].  Expected %x, got %x.", 6'd13, O[0][1][2]);
        end
        I[2][8][0] <= 6'd37;
        I[2][8][1] <= 6'd15;
        I[2][8][2] <= 6'd42;
        #1;
        if (!(O[2][8][0] === 6'd37)) begin
            $error("Failed on action=81 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][0].  Expected %x, got %x.", 6'd37, O[2][8][0]);
        end
        if (!(O[2][8][1] === 6'd15)) begin
            $error("Failed on action=82 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][1].  Expected %x, got %x.", 6'd15, O[2][8][1]);
        end
        if (!(O[2][8][2] === 6'd42)) begin
            $error("Failed on action=83 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][2].  Expected %x, got %x.", 6'd42, O[2][8][2]);
        end
        I[4][3][0] <= 6'd36;
        I[4][3][1] <= 6'd56;
        I[4][3][2] <= 6'd11;
        #1;
        if (!(O[4][3][0] === 6'd36)) begin
            $error("Failed on action=88 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][0].  Expected %x, got %x.", 6'd36, O[4][3][0]);
        end
        if (!(O[4][3][1] === 6'd56)) begin
            $error("Failed on action=89 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][1].  Expected %x, got %x.", 6'd56, O[4][3][1]);
        end
        if (!(O[4][3][2] === 6'd11)) begin
            $error("Failed on action=90 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][2].  Expected %x, got %x.", 6'd11, O[4][3][2]);
        end
        I[4][6][0] <= 6'd40;
        I[4][6][1] <= 6'd30;
        I[4][6][2] <= 6'd37;
        #1;
        if (!(O[4][6][0] === 6'd40)) begin
            $error("Failed on action=95 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][6][0].  Expected %x, got %x.", 6'd40, O[4][6][0]);
        end
        if (!(O[4][6][1] === 6'd30)) begin
            $error("Failed on action=96 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][6][1].  Expected %x, got %x.", 6'd30, O[4][6][1]);
        end
        if (!(O[4][6][2] === 6'd37)) begin
            $error("Failed on action=97 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][6][2].  Expected %x, got %x.", 6'd37, O[4][6][2]);
        end
        I[1][3][0] <= 6'd23;
        I[1][3][1] <= 6'd4;
        I[1][3][2] <= 6'd33;
        #1;
        if (!(O[1][3][0] === 6'd23)) begin
            $error("Failed on action=102 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][3][0].  Expected %x, got %x.", 6'd23, O[1][3][0]);
        end
        if (!(O[1][3][1] === 6'd4)) begin
            $error("Failed on action=103 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][3][1].  Expected %x, got %x.", 6'd4, O[1][3][1]);
        end
        if (!(O[1][3][2] === 6'd33)) begin
            $error("Failed on action=104 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][3][2].  Expected %x, got %x.", 6'd33, O[1][3][2]);
        end
        I[3][1][0] <= 6'd11;
        I[3][1][1] <= 6'd16;
        I[3][1][2] <= 6'd19;
        #1;
        if (!(O[3][1][0] === 6'd11)) begin
            $error("Failed on action=109 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][0].  Expected %x, got %x.", 6'd11, O[3][1][0]);
        end
        if (!(O[3][1][1] === 6'd16)) begin
            $error("Failed on action=110 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][1].  Expected %x, got %x.", 6'd16, O[3][1][1]);
        end
        if (!(O[3][1][2] === 6'd19)) begin
            $error("Failed on action=111 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][2].  Expected %x, got %x.", 6'd19, O[3][1][2]);
        end
        I[0][1][0] <= 6'd50;
        I[0][1][1] <= 6'd35;
        I[0][1][2] <= 6'd30;
        #1;
        if (!(O[0][1][0] === 6'd50)) begin
            $error("Failed on action=116 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][0].  Expected %x, got %x.", 6'd50, O[0][1][0]);
        end
        if (!(O[0][1][1] === 6'd35)) begin
            $error("Failed on action=117 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][1].  Expected %x, got %x.", 6'd35, O[0][1][1]);
        end
        if (!(O[0][1][2] === 6'd30)) begin
            $error("Failed on action=118 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][2].  Expected %x, got %x.", 6'd30, O[0][1][2]);
        end
        I[1][10][0] <= 6'd53;
        I[1][10][1] <= 6'd35;
        I[1][10][2] <= 6'd57;
        #1;
        if (!(O[1][10][0] === 6'd53)) begin
            $error("Failed on action=123 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][0].  Expected %x, got %x.", 6'd53, O[1][10][0]);
        end
        if (!(O[1][10][1] === 6'd35)) begin
            $error("Failed on action=124 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][1].  Expected %x, got %x.", 6'd35, O[1][10][1]);
        end
        if (!(O[1][10][2] === 6'd57)) begin
            $error("Failed on action=125 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][2].  Expected %x, got %x.", 6'd57, O[1][10][2]);
        end
        I[3][10][0] <= 6'd45;
        I[3][10][1] <= 6'd10;
        I[3][10][2] <= 6'd41;
        #1;
        if (!(O[3][10][0] === 6'd45)) begin
            $error("Failed on action=130 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][0].  Expected %x, got %x.", 6'd45, O[3][10][0]);
        end
        if (!(O[3][10][1] === 6'd10)) begin
            $error("Failed on action=131 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][1].  Expected %x, got %x.", 6'd10, O[3][10][1]);
        end
        if (!(O[3][10][2] === 6'd41)) begin
            $error("Failed on action=132 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][2].  Expected %x, got %x.", 6'd41, O[3][10][2]);
        end
        I[4][1][0] <= 6'd62;
        I[4][1][1] <= 6'd42;
        I[4][1][2] <= 6'd24;
        #1;
        if (!(O[4][1][0] === 6'd62)) begin
            $error("Failed on action=137 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][1][0].  Expected %x, got %x.", 6'd62, O[4][1][0]);
        end
        if (!(O[4][1][1] === 6'd42)) begin
            $error("Failed on action=138 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][1][1].  Expected %x, got %x.", 6'd42, O[4][1][1]);
        end
        if (!(O[4][1][2] === 6'd24)) begin
            $error("Failed on action=139 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][1][2].  Expected %x, got %x.", 6'd24, O[4][1][2]);
        end
        I[1][0][0] <= 6'd34;
        I[1][0][1] <= 6'd14;
        I[1][0][2] <= 6'd28;
        #1;
        if (!(O[1][0][0] === 6'd34)) begin
            $error("Failed on action=144 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][0].  Expected %x, got %x.", 6'd34, O[1][0][0]);
        end
        if (!(O[1][0][1] === 6'd14)) begin
            $error("Failed on action=145 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][1].  Expected %x, got %x.", 6'd14, O[1][0][1]);
        end
        if (!(O[1][0][2] === 6'd28)) begin
            $error("Failed on action=146 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][2].  Expected %x, got %x.", 6'd28, O[1][0][2]);
        end
        I[2][2][0] <= 6'd42;
        I[2][2][1] <= 6'd54;
        I[2][2][2] <= 6'd7;
        #1;
        if (!(O[2][2][0] === 6'd42)) begin
            $error("Failed on action=151 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][2][0].  Expected %x, got %x.", 6'd42, O[2][2][0]);
        end
        if (!(O[2][2][1] === 6'd54)) begin
            $error("Failed on action=152 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][2][1].  Expected %x, got %x.", 6'd54, O[2][2][1]);
        end
        if (!(O[2][2][2] === 6'd7)) begin
            $error("Failed on action=153 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][2][2].  Expected %x, got %x.", 6'd7, O[2][2][2]);
        end
        I[0][2][0] <= 6'd28;
        I[0][2][1] <= 6'd5;
        I[0][2][2] <= 6'd9;
        #1;
        if (!(O[0][2][0] === 6'd28)) begin
            $error("Failed on action=158 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][2][0].  Expected %x, got %x.", 6'd28, O[0][2][0]);
        end
        if (!(O[0][2][1] === 6'd5)) begin
            $error("Failed on action=159 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][2][1].  Expected %x, got %x.", 6'd5, O[0][2][1]);
        end
        if (!(O[0][2][2] === 6'd9)) begin
            $error("Failed on action=160 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][2][2].  Expected %x, got %x.", 6'd9, O[0][2][2]);
        end
        I[0][1][0] <= 6'd24;
        I[0][1][1] <= 6'd15;
        I[0][1][2] <= 6'd50;
        #1;
        if (!(O[0][1][0] === 6'd24)) begin
            $error("Failed on action=165 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][0].  Expected %x, got %x.", 6'd24, O[0][1][0]);
        end
        if (!(O[0][1][1] === 6'd15)) begin
            $error("Failed on action=166 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][1].  Expected %x, got %x.", 6'd15, O[0][1][1]);
        end
        if (!(O[0][1][2] === 6'd50)) begin
            $error("Failed on action=167 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][2].  Expected %x, got %x.", 6'd50, O[0][1][2]);
        end
        I[0][5][0] <= 6'd14;
        I[0][5][1] <= 6'd4;
        I[0][5][2] <= 6'd2;
        #1;
        if (!(O[0][5][0] === 6'd14)) begin
            $error("Failed on action=172 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][0].  Expected %x, got %x.", 6'd14, O[0][5][0]);
        end
        if (!(O[0][5][1] === 6'd4)) begin
            $error("Failed on action=173 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][1].  Expected %x, got %x.", 6'd4, O[0][5][1]);
        end
        if (!(O[0][5][2] === 6'd2)) begin
            $error("Failed on action=174 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][2].  Expected %x, got %x.", 6'd2, O[0][5][2]);
        end
        I[1][2][0] <= 6'd15;
        I[1][2][1] <= 6'd61;
        I[1][2][2] <= 6'd26;
        #1;
        if (!(O[1][2][0] === 6'd15)) begin
            $error("Failed on action=179 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][0].  Expected %x, got %x.", 6'd15, O[1][2][0]);
        end
        if (!(O[1][2][1] === 6'd61)) begin
            $error("Failed on action=180 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][1].  Expected %x, got %x.", 6'd61, O[1][2][1]);
        end
        if (!(O[1][2][2] === 6'd26)) begin
            $error("Failed on action=181 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][2].  Expected %x, got %x.", 6'd26, O[1][2][2]);
        end
        I[0][10][0] <= 6'd2;
        I[0][10][1] <= 6'd54;
        I[0][10][2] <= 6'd12;
        #1;
        if (!(O[0][10][0] === 6'd2)) begin
            $error("Failed on action=186 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][0].  Expected %x, got %x.", 6'd2, O[0][10][0]);
        end
        if (!(O[0][10][1] === 6'd54)) begin
            $error("Failed on action=187 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][1].  Expected %x, got %x.", 6'd54, O[0][10][1]);
        end
        if (!(O[0][10][2] === 6'd12)) begin
            $error("Failed on action=188 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][2].  Expected %x, got %x.", 6'd12, O[0][10][2]);
        end
        I[2][1][0] <= 6'd28;
        I[2][1][1] <= 6'd9;
        I[2][1][2] <= 6'd38;
        #1;
        if (!(O[2][1][0] === 6'd28)) begin
            $error("Failed on action=193 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][0].  Expected %x, got %x.", 6'd28, O[2][1][0]);
        end
        if (!(O[2][1][1] === 6'd9)) begin
            $error("Failed on action=194 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][1].  Expected %x, got %x.", 6'd9, O[2][1][1]);
        end
        if (!(O[2][1][2] === 6'd38)) begin
            $error("Failed on action=195 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][2].  Expected %x, got %x.", 6'd38, O[2][1][2]);
        end
        I[2][6][0] <= 6'd23;
        I[2][6][1] <= 6'd7;
        I[2][6][2] <= 6'd59;
        #1;
        if (!(O[2][6][0] === 6'd23)) begin
            $error("Failed on action=200 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][0].  Expected %x, got %x.", 6'd23, O[2][6][0]);
        end
        if (!(O[2][6][1] === 6'd7)) begin
            $error("Failed on action=201 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][1].  Expected %x, got %x.", 6'd7, O[2][6][1]);
        end
        if (!(O[2][6][2] === 6'd59)) begin
            $error("Failed on action=202 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][2].  Expected %x, got %x.", 6'd59, O[2][6][2]);
        end
        I[0][9][0] <= 6'd12;
        I[0][9][1] <= 6'd50;
        I[0][9][2] <= 6'd25;
        #1;
        if (!(O[0][9][0] === 6'd12)) begin
            $error("Failed on action=207 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][0].  Expected %x, got %x.", 6'd12, O[0][9][0]);
        end
        if (!(O[0][9][1] === 6'd50)) begin
            $error("Failed on action=208 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][1].  Expected %x, got %x.", 6'd50, O[0][9][1]);
        end
        if (!(O[0][9][2] === 6'd25)) begin
            $error("Failed on action=209 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][2].  Expected %x, got %x.", 6'd25, O[0][9][2]);
        end
        I[2][5][0] <= 6'd60;
        I[2][5][1] <= 6'd21;
        I[2][5][2] <= 6'd26;
        #1;
        if (!(O[2][5][0] === 6'd60)) begin
            $error("Failed on action=214 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][0].  Expected %x, got %x.", 6'd60, O[2][5][0]);
        end
        if (!(O[2][5][1] === 6'd21)) begin
            $error("Failed on action=215 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][1].  Expected %x, got %x.", 6'd21, O[2][5][1]);
        end
        if (!(O[2][5][2] === 6'd26)) begin
            $error("Failed on action=216 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][2].  Expected %x, got %x.", 6'd26, O[2][5][2]);
        end
        I[0][10][0] <= 6'd20;
        I[0][10][1] <= 6'd20;
        I[0][10][2] <= 6'd43;
        #1;
        if (!(O[0][10][0] === 6'd20)) begin
            $error("Failed on action=221 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][0].  Expected %x, got %x.", 6'd20, O[0][10][0]);
        end
        if (!(O[0][10][1] === 6'd20)) begin
            $error("Failed on action=222 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][1].  Expected %x, got %x.", 6'd20, O[0][10][1]);
        end
        if (!(O[0][10][2] === 6'd43)) begin
            $error("Failed on action=223 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][2].  Expected %x, got %x.", 6'd43, O[0][10][2]);
        end
        I[4][4][0] <= 6'd15;
        I[4][4][1] <= 6'd56;
        I[4][4][2] <= 6'd22;
        #1;
        if (!(O[4][4][0] === 6'd15)) begin
            $error("Failed on action=228 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][0].  Expected %x, got %x.", 6'd15, O[4][4][0]);
        end
        if (!(O[4][4][1] === 6'd56)) begin
            $error("Failed on action=229 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][1].  Expected %x, got %x.", 6'd56, O[4][4][1]);
        end
        if (!(O[4][4][2] === 6'd22)) begin
            $error("Failed on action=230 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][2].  Expected %x, got %x.", 6'd22, O[4][4][2]);
        end
        I[0][7][0] <= 6'd52;
        I[0][7][1] <= 6'd39;
        I[0][7][2] <= 6'd45;
        #1;
        if (!(O[0][7][0] === 6'd52)) begin
            $error("Failed on action=235 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][7][0].  Expected %x, got %x.", 6'd52, O[0][7][0]);
        end
        if (!(O[0][7][1] === 6'd39)) begin
            $error("Failed on action=236 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][7][1].  Expected %x, got %x.", 6'd39, O[0][7][1]);
        end
        if (!(O[0][7][2] === 6'd45)) begin
            $error("Failed on action=237 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][7][2].  Expected %x, got %x.", 6'd45, O[0][7][2]);
        end
        I[3][10][0] <= 6'd32;
        I[3][10][1] <= 6'd19;
        I[3][10][2] <= 6'd1;
        #1;
        if (!(O[3][10][0] === 6'd32)) begin
            $error("Failed on action=242 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][0].  Expected %x, got %x.", 6'd32, O[3][10][0]);
        end
        if (!(O[3][10][1] === 6'd19)) begin
            $error("Failed on action=243 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][1].  Expected %x, got %x.", 6'd19, O[3][10][1]);
        end
        if (!(O[3][10][2] === 6'd1)) begin
            $error("Failed on action=244 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][2].  Expected %x, got %x.", 6'd1, O[3][10][2]);
        end
        I[3][11][0] <= 6'd10;
        I[3][11][1] <= 6'd42;
        I[3][11][2] <= 6'd5;
        #1;
        if (!(O[3][11][0] === 6'd10)) begin
            $error("Failed on action=249 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][11][0].  Expected %x, got %x.", 6'd10, O[3][11][0]);
        end
        if (!(O[3][11][1] === 6'd42)) begin
            $error("Failed on action=250 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][11][1].  Expected %x, got %x.", 6'd42, O[3][11][1]);
        end
        if (!(O[3][11][2] === 6'd5)) begin
            $error("Failed on action=251 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][11][2].  Expected %x, got %x.", 6'd5, O[3][11][2]);
        end
        I[4][4][0] <= 6'd17;
        I[4][4][1] <= 6'd30;
        I[4][4][2] <= 6'd61;
        #1;
        if (!(O[4][4][0] === 6'd17)) begin
            $error("Failed on action=256 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][0].  Expected %x, got %x.", 6'd17, O[4][4][0]);
        end
        if (!(O[4][4][1] === 6'd30)) begin
            $error("Failed on action=257 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][1].  Expected %x, got %x.", 6'd30, O[4][4][1]);
        end
        if (!(O[4][4][2] === 6'd61)) begin
            $error("Failed on action=258 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][2].  Expected %x, got %x.", 6'd61, O[4][4][2]);
        end
        I[2][9][0] <= 6'd36;
        I[2][9][1] <= 6'd45;
        I[2][9][2] <= 6'd16;
        #1;
        if (!(O[2][9][0] === 6'd36)) begin
            $error("Failed on action=263 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][0].  Expected %x, got %x.", 6'd36, O[2][9][0]);
        end
        if (!(O[2][9][1] === 6'd45)) begin
            $error("Failed on action=264 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][1].  Expected %x, got %x.", 6'd45, O[2][9][1]);
        end
        if (!(O[2][9][2] === 6'd16)) begin
            $error("Failed on action=265 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][2].  Expected %x, got %x.", 6'd16, O[2][9][2]);
        end
        I[2][6][0] <= 6'd53;
        I[2][6][1] <= 6'd10;
        I[2][6][2] <= 6'd0;
        #1;
        if (!(O[2][6][0] === 6'd53)) begin
            $error("Failed on action=270 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][0].  Expected %x, got %x.", 6'd53, O[2][6][0]);
        end
        if (!(O[2][6][1] === 6'd10)) begin
            $error("Failed on action=271 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][1].  Expected %x, got %x.", 6'd10, O[2][6][1]);
        end
        if (!(O[2][6][2] === 6'd0)) begin
            $error("Failed on action=272 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][2].  Expected %x, got %x.", 6'd0, O[2][6][2]);
        end
        I[4][3][0] <= 6'd42;
        I[4][3][1] <= 6'd20;
        I[4][3][2] <= 6'd30;
        #1;
        if (!(O[4][3][0] === 6'd42)) begin
            $error("Failed on action=277 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][0].  Expected %x, got %x.", 6'd42, O[4][3][0]);
        end
        if (!(O[4][3][1] === 6'd20)) begin
            $error("Failed on action=278 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][1].  Expected %x, got %x.", 6'd20, O[4][3][1]);
        end
        if (!(O[4][3][2] === 6'd30)) begin
            $error("Failed on action=279 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][3][2].  Expected %x, got %x.", 6'd30, O[4][3][2]);
        end
        I[1][10][0] <= 6'd57;
        I[1][10][1] <= 6'd48;
        I[1][10][2] <= 6'd53;
        #1;
        if (!(O[1][10][0] === 6'd57)) begin
            $error("Failed on action=284 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][0].  Expected %x, got %x.", 6'd57, O[1][10][0]);
        end
        if (!(O[1][10][1] === 6'd48)) begin
            $error("Failed on action=285 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][1].  Expected %x, got %x.", 6'd48, O[1][10][1]);
        end
        if (!(O[1][10][2] === 6'd53)) begin
            $error("Failed on action=286 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][2].  Expected %x, got %x.", 6'd53, O[1][10][2]);
        end
        I[0][6][0] <= 6'd53;
        I[0][6][1] <= 6'd5;
        I[0][6][2] <= 6'd21;
        #1;
        if (!(O[0][6][0] === 6'd53)) begin
            $error("Failed on action=291 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][6][0].  Expected %x, got %x.", 6'd53, O[0][6][0]);
        end
        if (!(O[0][6][1] === 6'd5)) begin
            $error("Failed on action=292 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][6][1].  Expected %x, got %x.", 6'd5, O[0][6][1]);
        end
        if (!(O[0][6][2] === 6'd21)) begin
            $error("Failed on action=293 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][6][2].  Expected %x, got %x.", 6'd21, O[0][6][2]);
        end
        I[3][1][0] <= 6'd33;
        I[3][1][1] <= 6'd20;
        I[3][1][2] <= 6'd57;
        #1;
        if (!(O[3][1][0] === 6'd33)) begin
            $error("Failed on action=298 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][0].  Expected %x, got %x.", 6'd33, O[3][1][0]);
        end
        if (!(O[3][1][1] === 6'd20)) begin
            $error("Failed on action=299 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][1].  Expected %x, got %x.", 6'd20, O[3][1][1]);
        end
        if (!(O[3][1][2] === 6'd57)) begin
            $error("Failed on action=300 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][2].  Expected %x, got %x.", 6'd57, O[3][1][2]);
        end
        I[4][7][0] <= 6'd0;
        I[4][7][1] <= 6'd4;
        I[4][7][2] <= 6'd63;
        #1;
        if (!(O[4][7][0] === 6'd0)) begin
            $error("Failed on action=305 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][0].  Expected %x, got %x.", 6'd0, O[4][7][0]);
        end
        if (!(O[4][7][1] === 6'd4)) begin
            $error("Failed on action=306 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][1].  Expected %x, got %x.", 6'd4, O[4][7][1]);
        end
        if (!(O[4][7][2] === 6'd63)) begin
            $error("Failed on action=307 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][2].  Expected %x, got %x.", 6'd63, O[4][7][2]);
        end
        I[2][4][0] <= 6'd59;
        I[2][4][1] <= 6'd6;
        I[2][4][2] <= 6'd53;
        #1;
        if (!(O[2][4][0] === 6'd59)) begin
            $error("Failed on action=312 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][4][0].  Expected %x, got %x.", 6'd59, O[2][4][0]);
        end
        if (!(O[2][4][1] === 6'd6)) begin
            $error("Failed on action=313 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][4][1].  Expected %x, got %x.", 6'd6, O[2][4][1]);
        end
        if (!(O[2][4][2] === 6'd53)) begin
            $error("Failed on action=314 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][4][2].  Expected %x, got %x.", 6'd53, O[2][4][2]);
        end
        I[1][8][0] <= 6'd10;
        I[1][8][1] <= 6'd16;
        I[1][8][2] <= 6'd1;
        #1;
        if (!(O[1][8][0] === 6'd10)) begin
            $error("Failed on action=319 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][8][0].  Expected %x, got %x.", 6'd10, O[1][8][0]);
        end
        if (!(O[1][8][1] === 6'd16)) begin
            $error("Failed on action=320 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][8][1].  Expected %x, got %x.", 6'd16, O[1][8][1]);
        end
        if (!(O[1][8][2] === 6'd1)) begin
            $error("Failed on action=321 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][8][2].  Expected %x, got %x.", 6'd1, O[1][8][2]);
        end
        I[3][10][0] <= 6'd53;
        I[3][10][1] <= 6'd40;
        I[3][10][2] <= 6'd0;
        #1;
        if (!(O[3][10][0] === 6'd53)) begin
            $error("Failed on action=326 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][0].  Expected %x, got %x.", 6'd53, O[3][10][0]);
        end
        if (!(O[3][10][1] === 6'd40)) begin
            $error("Failed on action=327 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][1].  Expected %x, got %x.", 6'd40, O[3][10][1]);
        end
        if (!(O[3][10][2] === 6'd0)) begin
            $error("Failed on action=328 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][10][2].  Expected %x, got %x.", 6'd0, O[3][10][2]);
        end
        I[1][0][0] <= 6'd0;
        I[1][0][1] <= 6'd12;
        I[1][0][2] <= 6'd24;
        #1;
        if (!(O[1][0][0] === 6'd0)) begin
            $error("Failed on action=333 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][0].  Expected %x, got %x.", 6'd0, O[1][0][0]);
        end
        if (!(O[1][0][1] === 6'd12)) begin
            $error("Failed on action=334 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][1].  Expected %x, got %x.", 6'd12, O[1][0][1]);
        end
        if (!(O[1][0][2] === 6'd24)) begin
            $error("Failed on action=335 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][2].  Expected %x, got %x.", 6'd24, O[1][0][2]);
        end
        I[0][9][0] <= 6'd25;
        I[0][9][1] <= 6'd38;
        I[0][9][2] <= 6'd35;
        #1;
        if (!(O[0][9][0] === 6'd25)) begin
            $error("Failed on action=340 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][0].  Expected %x, got %x.", 6'd25, O[0][9][0]);
        end
        if (!(O[0][9][1] === 6'd38)) begin
            $error("Failed on action=341 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][1].  Expected %x, got %x.", 6'd38, O[0][9][1]);
        end
        if (!(O[0][9][2] === 6'd35)) begin
            $error("Failed on action=342 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][9][2].  Expected %x, got %x.", 6'd35, O[0][9][2]);
        end
        I[1][1][0] <= 6'd60;
        I[1][1][1] <= 6'd50;
        I[1][1][2] <= 6'd10;
        #1;
        if (!(O[1][1][0] === 6'd60)) begin
            $error("Failed on action=347 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][1][0].  Expected %x, got %x.", 6'd60, O[1][1][0]);
        end
        if (!(O[1][1][1] === 6'd50)) begin
            $error("Failed on action=348 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][1][1].  Expected %x, got %x.", 6'd50, O[1][1][1]);
        end
        if (!(O[1][1][2] === 6'd10)) begin
            $error("Failed on action=349 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][1][2].  Expected %x, got %x.", 6'd10, O[1][1][2]);
        end
        I[0][4][0] <= 6'd57;
        I[0][4][1] <= 6'd14;
        I[0][4][2] <= 6'd32;
        #1;
        if (!(O[0][4][0] === 6'd57)) begin
            $error("Failed on action=354 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][0].  Expected %x, got %x.", 6'd57, O[0][4][0]);
        end
        if (!(O[0][4][1] === 6'd14)) begin
            $error("Failed on action=355 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][1].  Expected %x, got %x.", 6'd14, O[0][4][1]);
        end
        if (!(O[0][4][2] === 6'd32)) begin
            $error("Failed on action=356 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][2].  Expected %x, got %x.", 6'd32, O[0][4][2]);
        end
        I[1][10][0] <= 6'd44;
        I[1][10][1] <= 6'd14;
        I[1][10][2] <= 6'd19;
        #1;
        if (!(O[1][10][0] === 6'd44)) begin
            $error("Failed on action=361 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][0].  Expected %x, got %x.", 6'd44, O[1][10][0]);
        end
        if (!(O[1][10][1] === 6'd14)) begin
            $error("Failed on action=362 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][1].  Expected %x, got %x.", 6'd14, O[1][10][1]);
        end
        if (!(O[1][10][2] === 6'd19)) begin
            $error("Failed on action=363 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][2].  Expected %x, got %x.", 6'd19, O[1][10][2]);
        end
        I[2][0][0] <= 6'd5;
        I[2][0][1] <= 6'd5;
        I[2][0][2] <= 6'd26;
        #1;
        if (!(O[2][0][0] === 6'd5)) begin
            $error("Failed on action=368 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][0][0].  Expected %x, got %x.", 6'd5, O[2][0][0]);
        end
        if (!(O[2][0][1] === 6'd5)) begin
            $error("Failed on action=369 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][0][1].  Expected %x, got %x.", 6'd5, O[2][0][1]);
        end
        if (!(O[2][0][2] === 6'd26)) begin
            $error("Failed on action=370 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][0][2].  Expected %x, got %x.", 6'd26, O[2][0][2]);
        end
        I[2][8][0] <= 6'd40;
        I[2][8][1] <= 6'd46;
        I[2][8][2] <= 6'd5;
        #1;
        if (!(O[2][8][0] === 6'd40)) begin
            $error("Failed on action=375 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][0].  Expected %x, got %x.", 6'd40, O[2][8][0]);
        end
        if (!(O[2][8][1] === 6'd46)) begin
            $error("Failed on action=376 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][1].  Expected %x, got %x.", 6'd46, O[2][8][1]);
        end
        if (!(O[2][8][2] === 6'd5)) begin
            $error("Failed on action=377 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][2].  Expected %x, got %x.", 6'd5, O[2][8][2]);
        end
        I[4][10][0] <= 6'd63;
        I[4][10][1] <= 6'd58;
        I[4][10][2] <= 6'd55;
        #1;
        if (!(O[4][10][0] === 6'd63)) begin
            $error("Failed on action=382 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][10][0].  Expected %x, got %x.", 6'd63, O[4][10][0]);
        end
        if (!(O[4][10][1] === 6'd58)) begin
            $error("Failed on action=383 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][10][1].  Expected %x, got %x.", 6'd58, O[4][10][1]);
        end
        if (!(O[4][10][2] === 6'd55)) begin
            $error("Failed on action=384 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][10][2].  Expected %x, got %x.", 6'd55, O[4][10][2]);
        end
        I[2][8][0] <= 6'd22;
        I[2][8][1] <= 6'd26;
        I[2][8][2] <= 6'd48;
        #1;
        if (!(O[2][8][0] === 6'd22)) begin
            $error("Failed on action=389 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][0].  Expected %x, got %x.", 6'd22, O[2][8][0]);
        end
        if (!(O[2][8][1] === 6'd26)) begin
            $error("Failed on action=390 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][1].  Expected %x, got %x.", 6'd26, O[2][8][1]);
        end
        if (!(O[2][8][2] === 6'd48)) begin
            $error("Failed on action=391 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][8][2].  Expected %x, got %x.", 6'd48, O[2][8][2]);
        end
        I[4][4][0] <= 6'd1;
        I[4][4][1] <= 6'd17;
        I[4][4][2] <= 6'd19;
        #1;
        if (!(O[4][4][0] === 6'd1)) begin
            $error("Failed on action=396 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][0].  Expected %x, got %x.", 6'd1, O[4][4][0]);
        end
        if (!(O[4][4][1] === 6'd17)) begin
            $error("Failed on action=397 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][1].  Expected %x, got %x.", 6'd17, O[4][4][1]);
        end
        if (!(O[4][4][2] === 6'd19)) begin
            $error("Failed on action=398 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][2].  Expected %x, got %x.", 6'd19, O[4][4][2]);
        end
        I[2][5][0] <= 6'd43;
        I[2][5][1] <= 6'd47;
        I[2][5][2] <= 6'd11;
        #1;
        if (!(O[2][5][0] === 6'd43)) begin
            $error("Failed on action=403 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][0].  Expected %x, got %x.", 6'd43, O[2][5][0]);
        end
        if (!(O[2][5][1] === 6'd47)) begin
            $error("Failed on action=404 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][1].  Expected %x, got %x.", 6'd47, O[2][5][1]);
        end
        if (!(O[2][5][2] === 6'd11)) begin
            $error("Failed on action=405 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][5][2].  Expected %x, got %x.", 6'd11, O[2][5][2]);
        end
        I[2][9][0] <= 6'd4;
        I[2][9][1] <= 6'd5;
        I[2][9][2] <= 6'd34;
        #1;
        if (!(O[2][9][0] === 6'd4)) begin
            $error("Failed on action=410 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][0].  Expected %x, got %x.", 6'd4, O[2][9][0]);
        end
        if (!(O[2][9][1] === 6'd5)) begin
            $error("Failed on action=411 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][1].  Expected %x, got %x.", 6'd5, O[2][9][1]);
        end
        if (!(O[2][9][2] === 6'd34)) begin
            $error("Failed on action=412 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][9][2].  Expected %x, got %x.", 6'd34, O[2][9][2]);
        end
        I[1][2][0] <= 6'd37;
        I[1][2][1] <= 6'd46;
        I[1][2][2] <= 6'd50;
        #1;
        if (!(O[1][2][0] === 6'd37)) begin
            $error("Failed on action=417 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][0].  Expected %x, got %x.", 6'd37, O[1][2][0]);
        end
        if (!(O[1][2][1] === 6'd46)) begin
            $error("Failed on action=418 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][1].  Expected %x, got %x.", 6'd46, O[1][2][1]);
        end
        if (!(O[1][2][2] === 6'd50)) begin
            $error("Failed on action=419 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][2].  Expected %x, got %x.", 6'd50, O[1][2][2]);
        end
        I[4][2][0] <= 6'd37;
        I[4][2][1] <= 6'd14;
        I[4][2][2] <= 6'd61;
        #1;
        if (!(O[4][2][0] === 6'd37)) begin
            $error("Failed on action=424 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][0].  Expected %x, got %x.", 6'd37, O[4][2][0]);
        end
        if (!(O[4][2][1] === 6'd14)) begin
            $error("Failed on action=425 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][1].  Expected %x, got %x.", 6'd14, O[4][2][1]);
        end
        if (!(O[4][2][2] === 6'd61)) begin
            $error("Failed on action=426 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][2].  Expected %x, got %x.", 6'd61, O[4][2][2]);
        end
        I[1][0][0] <= 6'd39;
        I[1][0][1] <= 6'd22;
        I[1][0][2] <= 6'd9;
        #1;
        if (!(O[1][0][0] === 6'd39)) begin
            $error("Failed on action=431 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][0].  Expected %x, got %x.", 6'd39, O[1][0][0]);
        end
        if (!(O[1][0][1] === 6'd22)) begin
            $error("Failed on action=432 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][1].  Expected %x, got %x.", 6'd22, O[1][0][1]);
        end
        if (!(O[1][0][2] === 6'd9)) begin
            $error("Failed on action=433 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][2].  Expected %x, got %x.", 6'd9, O[1][0][2]);
        end
        I[2][6][0] <= 6'd42;
        I[2][6][1] <= 6'd38;
        I[2][6][2] <= 6'd53;
        #1;
        if (!(O[2][6][0] === 6'd42)) begin
            $error("Failed on action=438 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][0].  Expected %x, got %x.", 6'd42, O[2][6][0]);
        end
        if (!(O[2][6][1] === 6'd38)) begin
            $error("Failed on action=439 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][1].  Expected %x, got %x.", 6'd38, O[2][6][1]);
        end
        if (!(O[2][6][2] === 6'd53)) begin
            $error("Failed on action=440 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][6][2].  Expected %x, got %x.", 6'd53, O[2][6][2]);
        end
        I[0][1][0] <= 6'd61;
        I[0][1][1] <= 6'd60;
        I[0][1][2] <= 6'd43;
        #1;
        if (!(O[0][1][0] === 6'd61)) begin
            $error("Failed on action=445 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][0].  Expected %x, got %x.", 6'd61, O[0][1][0]);
        end
        if (!(O[0][1][1] === 6'd60)) begin
            $error("Failed on action=446 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][1].  Expected %x, got %x.", 6'd60, O[0][1][1]);
        end
        if (!(O[0][1][2] === 6'd43)) begin
            $error("Failed on action=447 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][2].  Expected %x, got %x.", 6'd43, O[0][1][2]);
        end
        I[2][1][0] <= 6'd61;
        I[2][1][1] <= 6'd14;
        I[2][1][2] <= 6'd63;
        #1;
        if (!(O[2][1][0] === 6'd61)) begin
            $error("Failed on action=452 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][0].  Expected %x, got %x.", 6'd61, O[2][1][0]);
        end
        if (!(O[2][1][1] === 6'd14)) begin
            $error("Failed on action=453 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][1].  Expected %x, got %x.", 6'd14, O[2][1][1]);
        end
        if (!(O[2][1][2] === 6'd63)) begin
            $error("Failed on action=454 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][1][2].  Expected %x, got %x.", 6'd63, O[2][1][2]);
        end
        I[3][0][0] <= 6'd38;
        I[3][0][1] <= 6'd42;
        I[3][0][2] <= 6'd19;
        #1;
        if (!(O[3][0][0] === 6'd38)) begin
            $error("Failed on action=459 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][0].  Expected %x, got %x.", 6'd38, O[3][0][0]);
        end
        if (!(O[3][0][1] === 6'd42)) begin
            $error("Failed on action=460 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][1].  Expected %x, got %x.", 6'd42, O[3][0][1]);
        end
        if (!(O[3][0][2] === 6'd19)) begin
            $error("Failed on action=461 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][2].  Expected %x, got %x.", 6'd19, O[3][0][2]);
        end
        I[1][10][0] <= 6'd48;
        I[1][10][1] <= 6'd11;
        I[1][10][2] <= 6'd8;
        #1;
        if (!(O[1][10][0] === 6'd48)) begin
            $error("Failed on action=466 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][0].  Expected %x, got %x.", 6'd48, O[1][10][0]);
        end
        if (!(O[1][10][1] === 6'd11)) begin
            $error("Failed on action=467 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][1].  Expected %x, got %x.", 6'd11, O[1][10][1]);
        end
        if (!(O[1][10][2] === 6'd8)) begin
            $error("Failed on action=468 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][10][2].  Expected %x, got %x.", 6'd8, O[1][10][2]);
        end
        I[0][3][0] <= 6'd28;
        I[0][3][1] <= 6'd7;
        I[0][3][2] <= 6'd49;
        #1;
        if (!(O[0][3][0] === 6'd28)) begin
            $error("Failed on action=473 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][3][0].  Expected %x, got %x.", 6'd28, O[0][3][0]);
        end
        if (!(O[0][3][1] === 6'd7)) begin
            $error("Failed on action=474 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][3][1].  Expected %x, got %x.", 6'd7, O[0][3][1]);
        end
        if (!(O[0][3][2] === 6'd49)) begin
            $error("Failed on action=475 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][3][2].  Expected %x, got %x.", 6'd49, O[0][3][2]);
        end
        I[0][1][0] <= 6'd50;
        I[0][1][1] <= 6'd37;
        I[0][1][2] <= 6'd57;
        #1;
        if (!(O[0][1][0] === 6'd50)) begin
            $error("Failed on action=480 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][0].  Expected %x, got %x.", 6'd50, O[0][1][0]);
        end
        if (!(O[0][1][1] === 6'd37)) begin
            $error("Failed on action=481 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][1].  Expected %x, got %x.", 6'd37, O[0][1][1]);
        end
        if (!(O[0][1][2] === 6'd57)) begin
            $error("Failed on action=482 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][1][2].  Expected %x, got %x.", 6'd57, O[0][1][2]);
        end
        I[3][9][0] <= 6'd27;
        I[3][9][1] <= 6'd54;
        I[3][9][2] <= 6'd10;
        #1;
        if (!(O[3][9][0] === 6'd27)) begin
            $error("Failed on action=487 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][0].  Expected %x, got %x.", 6'd27, O[3][9][0]);
        end
        if (!(O[3][9][1] === 6'd54)) begin
            $error("Failed on action=488 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][1].  Expected %x, got %x.", 6'd54, O[3][9][1]);
        end
        if (!(O[3][9][2] === 6'd10)) begin
            $error("Failed on action=489 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][2].  Expected %x, got %x.", 6'd10, O[3][9][2]);
        end
        I[2][3][0] <= 6'd33;
        I[2][3][1] <= 6'd21;
        I[2][3][2] <= 6'd55;
        #1;
        if (!(O[2][3][0] === 6'd33)) begin
            $error("Failed on action=494 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][0].  Expected %x, got %x.", 6'd33, O[2][3][0]);
        end
        if (!(O[2][3][1] === 6'd21)) begin
            $error("Failed on action=495 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][1].  Expected %x, got %x.", 6'd21, O[2][3][1]);
        end
        if (!(O[2][3][2] === 6'd55)) begin
            $error("Failed on action=496 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][3][2].  Expected %x, got %x.", 6'd55, O[2][3][2]);
        end
        I[1][5][0] <= 6'd14;
        I[1][5][1] <= 6'd8;
        I[1][5][2] <= 6'd3;
        #1;
        if (!(O[1][5][0] === 6'd14)) begin
            $error("Failed on action=501 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][0].  Expected %x, got %x.", 6'd14, O[1][5][0]);
        end
        if (!(O[1][5][1] === 6'd8)) begin
            $error("Failed on action=502 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][1].  Expected %x, got %x.", 6'd8, O[1][5][1]);
        end
        if (!(O[1][5][2] === 6'd3)) begin
            $error("Failed on action=503 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][2].  Expected %x, got %x.", 6'd3, O[1][5][2]);
        end
        I[4][7][0] <= 6'd25;
        I[4][7][1] <= 6'd15;
        I[4][7][2] <= 6'd63;
        #1;
        if (!(O[4][7][0] === 6'd25)) begin
            $error("Failed on action=508 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][0].  Expected %x, got %x.", 6'd25, O[4][7][0]);
        end
        if (!(O[4][7][1] === 6'd15)) begin
            $error("Failed on action=509 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][1].  Expected %x, got %x.", 6'd15, O[4][7][1]);
        end
        if (!(O[4][7][2] === 6'd63)) begin
            $error("Failed on action=510 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][7][2].  Expected %x, got %x.", 6'd63, O[4][7][2]);
        end
        I[3][4][0] <= 6'd26;
        I[3][4][1] <= 6'd5;
        I[3][4][2] <= 6'd27;
        #1;
        if (!(O[3][4][0] === 6'd26)) begin
            $error("Failed on action=515 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][0].  Expected %x, got %x.", 6'd26, O[3][4][0]);
        end
        if (!(O[3][4][1] === 6'd5)) begin
            $error("Failed on action=516 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][1].  Expected %x, got %x.", 6'd5, O[3][4][1]);
        end
        if (!(O[3][4][2] === 6'd27)) begin
            $error("Failed on action=517 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][2].  Expected %x, got %x.", 6'd27, O[3][4][2]);
        end
        I[4][2][0] <= 6'd13;
        I[4][2][1] <= 6'd25;
        I[4][2][2] <= 6'd58;
        #1;
        if (!(O[4][2][0] === 6'd13)) begin
            $error("Failed on action=522 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][0].  Expected %x, got %x.", 6'd13, O[4][2][0]);
        end
        if (!(O[4][2][1] === 6'd25)) begin
            $error("Failed on action=523 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][1].  Expected %x, got %x.", 6'd25, O[4][2][1]);
        end
        if (!(O[4][2][2] === 6'd58)) begin
            $error("Failed on action=524 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][2].  Expected %x, got %x.", 6'd58, O[4][2][2]);
        end
        I[3][5][0] <= 6'd19;
        I[3][5][1] <= 6'd13;
        I[3][5][2] <= 6'd62;
        #1;
        if (!(O[3][5][0] === 6'd19)) begin
            $error("Failed on action=529 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][5][0].  Expected %x, got %x.", 6'd19, O[3][5][0]);
        end
        if (!(O[3][5][1] === 6'd13)) begin
            $error("Failed on action=530 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][5][1].  Expected %x, got %x.", 6'd13, O[3][5][1]);
        end
        if (!(O[3][5][2] === 6'd62)) begin
            $error("Failed on action=531 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][5][2].  Expected %x, got %x.", 6'd62, O[3][5][2]);
        end
        I[1][9][0] <= 6'd51;
        I[1][9][1] <= 6'd54;
        I[1][9][2] <= 6'd63;
        #1;
        if (!(O[1][9][0] === 6'd51)) begin
            $error("Failed on action=536 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][9][0].  Expected %x, got %x.", 6'd51, O[1][9][0]);
        end
        if (!(O[1][9][1] === 6'd54)) begin
            $error("Failed on action=537 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][9][1].  Expected %x, got %x.", 6'd54, O[1][9][1]);
        end
        if (!(O[1][9][2] === 6'd63)) begin
            $error("Failed on action=538 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][9][2].  Expected %x, got %x.", 6'd63, O[1][9][2]);
        end
        I[2][7][0] <= 6'd63;
        I[2][7][1] <= 6'd25;
        I[2][7][2] <= 6'd28;
        #1;
        if (!(O[2][7][0] === 6'd63)) begin
            $error("Failed on action=543 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][7][0].  Expected %x, got %x.", 6'd63, O[2][7][0]);
        end
        if (!(O[2][7][1] === 6'd25)) begin
            $error("Failed on action=544 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][7][1].  Expected %x, got %x.", 6'd25, O[2][7][1]);
        end
        if (!(O[2][7][2] === 6'd28)) begin
            $error("Failed on action=545 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][7][2].  Expected %x, got %x.", 6'd28, O[2][7][2]);
        end
        I[0][5][0] <= 6'd40;
        I[0][5][1] <= 6'd41;
        I[0][5][2] <= 6'd4;
        #1;
        if (!(O[0][5][0] === 6'd40)) begin
            $error("Failed on action=550 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][0].  Expected %x, got %x.", 6'd40, O[0][5][0]);
        end
        if (!(O[0][5][1] === 6'd41)) begin
            $error("Failed on action=551 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][1].  Expected %x, got %x.", 6'd41, O[0][5][1]);
        end
        if (!(O[0][5][2] === 6'd4)) begin
            $error("Failed on action=552 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][5][2].  Expected %x, got %x.", 6'd4, O[0][5][2]);
        end
        I[4][2][0] <= 6'd32;
        I[4][2][1] <= 6'd19;
        I[4][2][2] <= 6'd48;
        #1;
        if (!(O[4][2][0] === 6'd32)) begin
            $error("Failed on action=557 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][0].  Expected %x, got %x.", 6'd32, O[4][2][0]);
        end
        if (!(O[4][2][1] === 6'd19)) begin
            $error("Failed on action=558 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][1].  Expected %x, got %x.", 6'd19, O[4][2][1]);
        end
        if (!(O[4][2][2] === 6'd48)) begin
            $error("Failed on action=559 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][2][2].  Expected %x, got %x.", 6'd48, O[4][2][2]);
        end
        I[4][4][0] <= 6'd60;
        I[4][4][1] <= 6'd8;
        I[4][4][2] <= 6'd10;
        #1;
        if (!(O[4][4][0] === 6'd60)) begin
            $error("Failed on action=564 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][0].  Expected %x, got %x.", 6'd60, O[4][4][0]);
        end
        if (!(O[4][4][1] === 6'd8)) begin
            $error("Failed on action=565 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][1].  Expected %x, got %x.", 6'd8, O[4][4][1]);
        end
        if (!(O[4][4][2] === 6'd10)) begin
            $error("Failed on action=566 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][4][2].  Expected %x, got %x.", 6'd10, O[4][4][2]);
        end
        I[4][0][0] <= 6'd8;
        I[4][0][1] <= 6'd28;
        I[4][0][2] <= 6'd16;
        #1;
        if (!(O[4][0][0] === 6'd8)) begin
            $error("Failed on action=571 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][0][0].  Expected %x, got %x.", 6'd8, O[4][0][0]);
        end
        if (!(O[4][0][1] === 6'd28)) begin
            $error("Failed on action=572 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][0][1].  Expected %x, got %x.", 6'd28, O[4][0][1]);
        end
        if (!(O[4][0][2] === 6'd16)) begin
            $error("Failed on action=573 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][0][2].  Expected %x, got %x.", 6'd16, O[4][0][2]);
        end
        I[0][4][0] <= 6'd1;
        I[0][4][1] <= 6'd57;
        I[0][4][2] <= 6'd42;
        #1;
        if (!(O[0][4][0] === 6'd1)) begin
            $error("Failed on action=578 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][0].  Expected %x, got %x.", 6'd1, O[0][4][0]);
        end
        if (!(O[0][4][1] === 6'd57)) begin
            $error("Failed on action=579 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][1].  Expected %x, got %x.", 6'd57, O[0][4][1]);
        end
        if (!(O[0][4][2] === 6'd42)) begin
            $error("Failed on action=580 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][4][2].  Expected %x, got %x.", 6'd42, O[0][4][2]);
        end
        I[1][2][0] <= 6'd58;
        I[1][2][1] <= 6'd47;
        I[1][2][2] <= 6'd48;
        #1;
        if (!(O[1][2][0] === 6'd58)) begin
            $error("Failed on action=585 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][0].  Expected %x, got %x.", 6'd58, O[1][2][0]);
        end
        if (!(O[1][2][1] === 6'd47)) begin
            $error("Failed on action=586 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][1].  Expected %x, got %x.", 6'd47, O[1][2][1]);
        end
        if (!(O[1][2][2] === 6'd48)) begin
            $error("Failed on action=587 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][2][2].  Expected %x, got %x.", 6'd48, O[1][2][2]);
        end
        I[4][8][0] <= 6'd4;
        I[4][8][1] <= 6'd11;
        I[4][8][2] <= 6'd9;
        #1;
        if (!(O[4][8][0] === 6'd4)) begin
            $error("Failed on action=592 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][8][0].  Expected %x, got %x.", 6'd4, O[4][8][0]);
        end
        if (!(O[4][8][1] === 6'd11)) begin
            $error("Failed on action=593 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][8][1].  Expected %x, got %x.", 6'd11, O[4][8][1]);
        end
        if (!(O[4][8][2] === 6'd9)) begin
            $error("Failed on action=594 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[4][8][2].  Expected %x, got %x.", 6'd9, O[4][8][2]);
        end
        I[3][3][0] <= 6'd37;
        I[3][3][1] <= 6'd53;
        I[3][3][2] <= 6'd61;
        #1;
        if (!(O[3][3][0] === 6'd37)) begin
            $error("Failed on action=599 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][3][0].  Expected %x, got %x.", 6'd37, O[3][3][0]);
        end
        if (!(O[3][3][1] === 6'd53)) begin
            $error("Failed on action=600 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][3][1].  Expected %x, got %x.", 6'd53, O[3][3][1]);
        end
        if (!(O[3][3][2] === 6'd61)) begin
            $error("Failed on action=601 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][3][2].  Expected %x, got %x.", 6'd61, O[3][3][2]);
        end
        I[3][9][0] <= 6'd29;
        I[3][9][1] <= 6'd2;
        I[3][9][2] <= 6'd0;
        #1;
        if (!(O[3][9][0] === 6'd29)) begin
            $error("Failed on action=606 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][0].  Expected %x, got %x.", 6'd29, O[3][9][0]);
        end
        if (!(O[3][9][1] === 6'd2)) begin
            $error("Failed on action=607 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][1].  Expected %x, got %x.", 6'd2, O[3][9][1]);
        end
        if (!(O[3][9][2] === 6'd0)) begin
            $error("Failed on action=608 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][9][2].  Expected %x, got %x.", 6'd0, O[3][9][2]);
        end
        I[1][4][0] <= 6'd32;
        I[1][4][1] <= 6'd42;
        I[1][4][2] <= 6'd8;
        #1;
        if (!(O[1][4][0] === 6'd32)) begin
            $error("Failed on action=613 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][4][0].  Expected %x, got %x.", 6'd32, O[1][4][0]);
        end
        if (!(O[1][4][1] === 6'd42)) begin
            $error("Failed on action=614 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][4][1].  Expected %x, got %x.", 6'd42, O[1][4][1]);
        end
        if (!(O[1][4][2] === 6'd8)) begin
            $error("Failed on action=615 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][4][2].  Expected %x, got %x.", 6'd8, O[1][4][2]);
        end
        I[3][4][0] <= 6'd38;
        I[3][4][1] <= 6'd52;
        I[3][4][2] <= 6'd49;
        #1;
        if (!(O[3][4][0] === 6'd38)) begin
            $error("Failed on action=620 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][0].  Expected %x, got %x.", 6'd38, O[3][4][0]);
        end
        if (!(O[3][4][1] === 6'd52)) begin
            $error("Failed on action=621 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][1].  Expected %x, got %x.", 6'd52, O[3][4][1]);
        end
        if (!(O[3][4][2] === 6'd49)) begin
            $error("Failed on action=622 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][4][2].  Expected %x, got %x.", 6'd49, O[3][4][2]);
        end
        I[3][0][0] <= 6'd20;
        I[3][0][1] <= 6'd16;
        I[3][0][2] <= 6'd30;
        #1;
        if (!(O[3][0][0] === 6'd20)) begin
            $error("Failed on action=627 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][0].  Expected %x, got %x.", 6'd20, O[3][0][0]);
        end
        if (!(O[3][0][1] === 6'd16)) begin
            $error("Failed on action=628 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][1].  Expected %x, got %x.", 6'd16, O[3][0][1]);
        end
        if (!(O[3][0][2] === 6'd30)) begin
            $error("Failed on action=629 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][0][2].  Expected %x, got %x.", 6'd30, O[3][0][2]);
        end
        I[2][11][0] <= 6'd42;
        I[2][11][1] <= 6'd7;
        I[2][11][2] <= 6'd4;
        #1;
        if (!(O[2][11][0] === 6'd42)) begin
            $error("Failed on action=634 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][0].  Expected %x, got %x.", 6'd42, O[2][11][0]);
        end
        if (!(O[2][11][1] === 6'd7)) begin
            $error("Failed on action=635 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][1].  Expected %x, got %x.", 6'd7, O[2][11][1]);
        end
        if (!(O[2][11][2] === 6'd4)) begin
            $error("Failed on action=636 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][2].  Expected %x, got %x.", 6'd4, O[2][11][2]);
        end
        I[3][6][0] <= 6'd18;
        I[3][6][1] <= 6'd62;
        I[3][6][2] <= 6'd10;
        #1;
        if (!(O[3][6][0] === 6'd18)) begin
            $error("Failed on action=641 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][0].  Expected %x, got %x.", 6'd18, O[3][6][0]);
        end
        if (!(O[3][6][1] === 6'd62)) begin
            $error("Failed on action=642 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][1].  Expected %x, got %x.", 6'd62, O[3][6][1]);
        end
        if (!(O[3][6][2] === 6'd10)) begin
            $error("Failed on action=643 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][6][2].  Expected %x, got %x.", 6'd10, O[3][6][2]);
        end
        I[1][5][0] <= 6'd52;
        I[1][5][1] <= 6'd4;
        I[1][5][2] <= 6'd59;
        #1;
        if (!(O[1][5][0] === 6'd52)) begin
            $error("Failed on action=648 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][0].  Expected %x, got %x.", 6'd52, O[1][5][0]);
        end
        if (!(O[1][5][1] === 6'd4)) begin
            $error("Failed on action=649 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][1].  Expected %x, got %x.", 6'd4, O[1][5][1]);
        end
        if (!(O[1][5][2] === 6'd59)) begin
            $error("Failed on action=650 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][5][2].  Expected %x, got %x.", 6'd59, O[1][5][2]);
        end
        I[3][7][0] <= 6'd6;
        I[3][7][1] <= 6'd12;
        I[3][7][2] <= 6'd60;
        #1;
        if (!(O[3][7][0] === 6'd6)) begin
            $error("Failed on action=655 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][0].  Expected %x, got %x.", 6'd6, O[3][7][0]);
        end
        if (!(O[3][7][1] === 6'd12)) begin
            $error("Failed on action=656 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][1].  Expected %x, got %x.", 6'd12, O[3][7][1]);
        end
        if (!(O[3][7][2] === 6'd60)) begin
            $error("Failed on action=657 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][2].  Expected %x, got %x.", 6'd60, O[3][7][2]);
        end
        I[1][0][0] <= 6'd4;
        I[1][0][1] <= 6'd16;
        I[1][0][2] <= 6'd41;
        #1;
        if (!(O[1][0][0] === 6'd4)) begin
            $error("Failed on action=662 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][0].  Expected %x, got %x.", 6'd4, O[1][0][0]);
        end
        if (!(O[1][0][1] === 6'd16)) begin
            $error("Failed on action=663 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][1].  Expected %x, got %x.", 6'd16, O[1][0][1]);
        end
        if (!(O[1][0][2] === 6'd41)) begin
            $error("Failed on action=664 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[1][0][2].  Expected %x, got %x.", 6'd41, O[1][0][2]);
        end
        I[0][11][0] <= 6'd44;
        I[0][11][1] <= 6'd24;
        I[0][11][2] <= 6'd49;
        #1;
        if (!(O[0][11][0] === 6'd44)) begin
            $error("Failed on action=669 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][0].  Expected %x, got %x.", 6'd44, O[0][11][0]);
        end
        if (!(O[0][11][1] === 6'd24)) begin
            $error("Failed on action=670 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][1].  Expected %x, got %x.", 6'd24, O[0][11][1]);
        end
        if (!(O[0][11][2] === 6'd49)) begin
            $error("Failed on action=671 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][11][2].  Expected %x, got %x.", 6'd49, O[0][11][2]);
        end
        I[3][1][0] <= 6'd7;
        I[3][1][1] <= 6'd59;
        I[3][1][2] <= 6'd43;
        #1;
        if (!(O[3][1][0] === 6'd7)) begin
            $error("Failed on action=676 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][0].  Expected %x, got %x.", 6'd7, O[3][1][0]);
        end
        if (!(O[3][1][1] === 6'd59)) begin
            $error("Failed on action=677 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][1].  Expected %x, got %x.", 6'd59, O[3][1][1]);
        end
        if (!(O[3][1][2] === 6'd43)) begin
            $error("Failed on action=678 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][1][2].  Expected %x, got %x.", 6'd43, O[3][1][2]);
        end
        I[0][10][0] <= 6'd37;
        I[0][10][1] <= 6'd16;
        I[0][10][2] <= 6'd49;
        #1;
        if (!(O[0][10][0] === 6'd37)) begin
            $error("Failed on action=683 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][0].  Expected %x, got %x.", 6'd37, O[0][10][0]);
        end
        if (!(O[0][10][1] === 6'd16)) begin
            $error("Failed on action=684 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][1].  Expected %x, got %x.", 6'd16, O[0][10][1]);
        end
        if (!(O[0][10][2] === 6'd49)) begin
            $error("Failed on action=685 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[0][10][2].  Expected %x, got %x.", 6'd49, O[0][10][2]);
        end
        I[2][11][0] <= 6'd15;
        I[2][11][1] <= 6'd24;
        I[2][11][2] <= 6'd4;
        #1;
        if (!(O[2][11][0] === 6'd15)) begin
            $error("Failed on action=690 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][0].  Expected %x, got %x.", 6'd15, O[2][11][0]);
        end
        if (!(O[2][11][1] === 6'd24)) begin
            $error("Failed on action=691 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][1].  Expected %x, got %x.", 6'd24, O[2][11][1]);
        end
        if (!(O[2][11][2] === 6'd4)) begin
            $error("Failed on action=692 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[2][11][2].  Expected %x, got %x.", 6'd4, O[2][11][2]);
        end
        I[3][7][0] <= 6'd47;
        I[3][7][1] <= 6'd24;
        I[3][7][2] <= 6'd58;
        #1;
        if (!(O[3][7][0] === 6'd47)) begin
            $error("Failed on action=697 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][0].  Expected %x, got %x.", 6'd47, O[3][7][0]);
        end
        if (!(O[3][7][1] === 6'd24)) begin
            $error("Failed on action=698 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][1].  Expected %x, got %x.", 6'd24, O[3][7][1]);
        end
        if (!(O[3][7][2] === 6'd58)) begin
            $error("Failed on action=699 checking port test_system_verilog_target_packed_arrays_False__test_packed_arrays_stimulate_bulk.O[3][7][2].  Expected %x, got %x.", 6'd58, O[3][7][2]);
        end

        #20 $finish;
    end

endmodule
