module error_task;
    initial begin
        $error;
        $finish;
    end
endmodule
