module mybuf(
    input in_,
    output out
);

    assign out = in_;

endmodule
