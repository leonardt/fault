module bidir(
    inout a,
    inout b
);

    tran tran_i(a, b);

endmodule
